parameter DIN_WIDTH=22;
parameter M=1;
parameter N=4;
parameter R=160;
parameter DOUT_WIDTH=54;
parameter MODE=0;

parameter DIN_WIDTH=18;
parameter M=1;
parameter N=5;
parameter R=16;
parameter DOUT_WIDTH=38;
parameter MODE=0;

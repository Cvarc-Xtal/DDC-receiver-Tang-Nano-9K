`define MODULE_NAME CIC_Filter_2
`define DECIMATOR

parameter DIN_WIDTH=24;
parameter M=1;
parameter N=4;
parameter R=2;
parameter DOUT_WIDTH=28;
parameter MODE=0;

`define MODULE_NAME CIC_Filter_d16
`define DECIMATOR

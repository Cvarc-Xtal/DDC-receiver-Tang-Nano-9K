`define MODULE_NAME CIC_Fliter_160
`define DECIMATOR
